library verilog;
use verilog.vl_types.all;
entity latch_32bit_vlg_vec_tst is
end latch_32bit_vlg_vec_tst;
