library verilog;
use verilog.vl_types.all;
entity mux_4to1_vlg_vec_tst is
end mux_4to1_vlg_vec_tst;
