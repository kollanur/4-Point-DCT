library verilog;
use verilog.vl_types.all;
entity adder_32bit_vlg_vec_tst is
end adder_32bit_vlg_vec_tst;
