library verilog;
use verilog.vl_types.all;
entity demux_1to2_vlg_vec_tst is
end demux_1to2_vlg_vec_tst;
