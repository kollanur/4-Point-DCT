library verilog;
use verilog.vl_types.all;
entity multiplier_32bit_vlg_vec_tst is
end multiplier_32bit_vlg_vec_tst;
